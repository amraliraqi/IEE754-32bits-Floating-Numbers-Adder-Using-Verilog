`timescale 1ns/1ps
module TB_NormalNumbers();

parameter DELAY=10;
reg [31:0] NumberA;
reg [31:0] NumberB;
reg A_S;  // zero for add, one for subb
wire [31:0] Result;

Final Final(NumberA,NumberB,A_S,Result);
initial
    begin
     
    // Normal Case 1:  (1.417843161699894*10^38) - (1.417842756051702*10^38) = 4.056481920730334*10^31
    NumberA = 32'b0_11111101_10101010101010101010101;
    NumberB = 32'b0_11111101_10101010101010101010001;
    A_S = 1'b1;
    #DELAY;

    if(Result == 32'b0_11101000_00000000000000000000000 )
            $display("Normal Case 1 passed     ,result is 4.056481920730334*10^31 = %b",Result);
    else
            $display("Normal Case 1 failed     ,result is 4.056481920730334*10^31 = %b",32'b0_11101000_00000000000000000000000);
             
    /*********************************************************************************************************/
    #DELAY;

    // Normal Case 2:  (4.422139697774293*10^35) - (5.538449850390212*10^35) = -1.116310152615919*10^35
    NumberA = 32'b0_11110101_01010100101010110101010;
    NumberB = 32'b0_11110101_10101010101010101010101;
    A_S = 1'b1;
    #DELAY;

    if(Result == 32'b1_11110011_01010111111111010101100 )
            $display("Normal Case 2 passed     ,result is -1.116310152615919*10^35 = %b",Result);
    else
            $display("Normal Case 2 failed     ,result is -1.116310152615919*10^35 = %b",32'b1_11110101_01010111111111010101100);
             
    /*********************************************************************************************************/
    #DELAY;

    // Normal Case 3:  (-1.701411733192644*10^37) + (1.415084703287774*10^37) = -2.863270299048707*10^36
    NumberA = 32'b1_11111010_10011001100110011001100;
    NumberB = 32'b0_11111010_01010100101010110101010;
    A_S = 1'b0;
    #DELAY;

    if(Result == 32'b1_11111000_00010011101110010001000 )
            $display("Normal Case 3 passed     ,result is -2.863270299048707*10^36 = %b",Result);
    else
            $display("Normal Case 3 failed     ,result is -2.863270299048707*10^36 = %b",32'b1_11111000_00010011101110010001000);

    /*********************************************************************************************************/
    #DELAY;

    // Normal Case 4:  (-1.799996137003937*10^34) + (-1.791851358103467*10^34) = -3.591847495107403*10^34
    NumberA = 32'b1_11110000_10111011101110111011101;
    NumberB = 32'b1_11110000_10111001101110011011100;
    A_S = 1'b0;
    #DELAY;

    if(Result == 32'b1_11110001_01110101011101010111001 )
            $display("Normal Case 4 passed     ,result is -3.591847495107403*10^34 =%b",Result);
    else
            $display("Normal Case 4 failed     ,result is -3.591847495107403*10^34 =%b",32'b1_11110001_01110101011101010111001);  

    /*********************************************************************************************************/
    #DELAY;
          

    $stop;
    end

endmodule

